`include "../Arithmetic.v"

module ADD16_tb;

    reg [15:0] A, B;
    wire [15:0]sum;

    ADD16 add16(.sum(sum), .A(A), .B(B));

    initial begin
            A = 16'b0000000000000000; B = 16'b0000000000000000; // out -> 0000000000000000
        #1  A = 16'b0000000000000000; B = 16'b1111111111111111; // out -> 1111111111111111
        #1  A = 16'b1111111111111111; B = 16'b1111111111111111; // out -> 1111111111111110
        #1  A = 16'b1010101010101010; B = 16'b0101010101010101; // out -> 1111111111111111
        #1  A = 16'b0011110011000011; B = 16'b0000111111110000; // out -> 0100110010110011
        #1  A = 16'b0001001000110100; B = 16'b1001100001110110; // out -> 1010101010101010
    end

    initial begin
        $monitor ("%t | A = %b | B = %b | sum = %b", $time, A, B, sum);
        $dumpfile("./DumpFiles/add16_dump.vcd");
        $dumpvars();
    end

endmodule